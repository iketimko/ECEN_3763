
module KEY (
	probe,
	source);	

	input	[3:0]	probe;
	output	[3:0]	source;
endmodule
