// KEY.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module KEY (
		input  wire [3:0] probe,  //  probes.probe
		output wire [3:0] source  // sources.source
	);

	altsource_probe_top #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("NONE"),
		.probe_width             (4),
		.source_width            (4),
		.source_initial_value    ("F"),
		.enable_metastability    ("NO")
	) in_system_sources_probes_0 (
		.source     (source), // sources.source
		.probe      (probe),  //  probes.probe
		.source_ena (1'b1)    // (terminated)
	);

endmodule
