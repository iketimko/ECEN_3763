//`ifdef _720p_resolution
    parameter HFP_WIDTH = 'd110;
    parameter HSYNCH_WIDTH = 'd40;
    parameter HBP_WIDTH = 'd220;
    parameter IMAGE_WIDTH = 'd1280;
    parameter VFP_HEIGHT = 'd5;
    parameter VSYNCH_HEIGHT = 'd5;
    parameter VBP_HEIGHT = 'd20;
    parameter IMAGE_HEIGHT = 'd720;
//`endif _720p_resolution

// `ifdef _1080p_resolution
    
// `endif _1080p_resolution