// PD_L12.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module PD_L12 (
		input  wire  clk_clk,             //           clk.clk
		output wire  pll_0_locked_export, //  pll_0_locked.export
		output wire  pll_0_outclk0_clk,   // pll_0_outclk0.clk
		input  wire  reset_reset_n        //         reset.reset_n
	);

	PD_L12_pll_0 pll_0 (
		.refclk   (clk_clk),             //  refclk.clk
		.rst      (~reset_reset_n),      //   reset.reset
		.outclk_0 (pll_0_outclk0_clk),   // outclk0.clk
		.locked   (pll_0_locked_export)  //  locked.export
	);

endmodule
