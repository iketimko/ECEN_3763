
module ISSP_IT_LAB_3 (
	source,
	probe);	

	output	[0:0]	source;
	input	[0:0]	probe;
endmodule
