module Test (input [0:0] KEY, output [0:0] LEDR);

assign LEDR[0] = KEY[0];

endmodule